* ON SEMICONDUCTOR NEXT GEN MODEL, JAN 2019
* BEGIN MODEL NCS2007
*
* MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT
* THROUGH THE SUPPLY RAILS, RAIL-TO-RAIL OUTPUT STAGE,
* OUTPUT CURRENT LIMIT, UNSYMETRICAL SLEW RATE WITH
* TEMPERATURE EFFECTS , OUTPUT SWING VERSUS CURRENT
* AND TEMPERATURE, OPEN LOOP GAIN AND PHASE WITH RL
* AND CL EFFECTS, POWER SUPPLY REJECTION WITH
* FREQUENCY EFFECTS, COMMON MODE REJECTION WITH
* FREQUENCY AND SUPPLY VOLTAGE EFFECTS, ROUGH SETTLING
* TIME, INPUT VOLTAGE NOISE, INPUT CURRENT NOISE,
* INPUT BIAS CURRENT WITH TEMPERATURE EFFECTS, INPUT
* CAPACITANCE, INPUT COMMON MODE RANGE, OFFSET WITH
* TEMPERATURE EFFECTS, INPUT AND OUTPUT CLAMPS TO
* THE RAILS, INPUT DIFFERENTIAL CLAMP, INPUT EMI
* FILTER, AND QUIESCENT CURRENT WITH VOLTAGE AND
* TEMPERATURE EFFECTS.
*
* MODEL TOTAL SUPPLY VOLTAGE RANGE IS 2.7 TO 36 V.
* MODEL TEMP RANGE IS -40 TO +125 DEG C.
* NOTE THAT MODEL IS FUNCTIONAL OVER THIS RANGE BUT
* NOT ALL PARAMETERS TRACK THOSE OF THE REAL PART.

* NOTE - FOR ACCURATE BIAS CURRENTS AT ROOM AND COLD
* SET THE SPICE ANALYSIS OPTIONS AS FOLLOWS:
* GMIN 1E-13, ABSTOL 1E-14, RELTOL 1E-6.
* ALL OF THESE OPTIONS ARE SMALLER THAN THE
* DEFAULTS IN MOST SIMULATORS, SET THEM ALL AS SMALL
* AS WILL ALLOW CONVERGANCE ON YOUR SIMULATOR.

* IF YOU ARE USING LTSPICE17 ADD THE OPTIONS
* PLOTRELTOL=1E-4 AND PLOTVNTOL=1E-6 FOR MORE
* ACCURATE TIME DOMAIN WAVEFORM PLOTTING.
*
* PINOUT  1    2    3    4    5
* PINOUT +IN  -IN  +V   -V   OUT
*
.SUBCKT NCS2007 1 2 3 4 5
Q20 195 196 112 QN
R3 197 198 2
R4 199 198 2
R10 196 200 1E3
R11 201 202 1E3
R12 203 3 0.335
R13 4 204 0.258
R17 205 110 0.335
R18 112 206 0.258
D7 207 0 DIN
D8 208 0 DIN
I8 0 207 12E-6
I9 0 208 12E-6
E2 112 0 4 0 1
E3 110 0 3 0 1
E4 209 2 210 211 0.068
G2 212 2 213 214 5.023E-7
E5 215 0 110 0 1
E6 216 0 112 0 1
E7 217 0 VCM 115 1
R30 215 218 1E6
R31 216 219 1E6
R32 217 220 1E6
R33 0 218 10
R34 0 219 10
R35 0 220 10
E10 144 221 220 0 4E-4
R36 222 VCM 1E3
R37 VCM 223 1E3
C6 215 218 15E-9
C7 216 219 15E-9
C8 217 220 400E-12
E11 224 1 219 0 -0.05
E12 212 224 218 0 0.05
E14 115 112 110 112 0.5
M1 225 113 204 204 NOUT L=3U W=1400U
M2 226 227 203 203 POUT L=3U W=1400U
M3 118 118 205 205 POUT L=3U W=1400U
M4 228 229 197 197 HVP L=30U W=6000U
M5 230 231 199 199 HVP L=30U W=6000U
M8 119 119 206 206 NOUT L=3U W=1400U
R43 111 227 300
R44 232 113 300
G3 114 115 233 115 3.33E-4
R45 115 114 1.2E9
R46 112 228 490
R47 112 230 490
C13 228 230 4.0E-12
C14 229 0 1.65E-12
C15 231 0 1.65E-12
C16 120 0 0.1E-12
D13 113 195 DB
D14 234 227 DB
Q15 234 201 110 QP
V18 235 229 1.37E-3
M19 236 237 238 238 PIN L=60U W=5000U
E17 223 0 212 0 1
E18 222 0 2 0 1
M23 237 237 238 238 PIN L=60U W=5000U
V21 236 239 0
R59 120 226 35 TC=3.48E-3,1.45E-5
R60 225 120 28 TC=3.48E-3,1.45E-5
J1 240 212 240 JC
J2 240 209 240 JC
J3 209 241 209 JC
J4 212 241 212 JC
C21 229 231 0.63E-12
E20 144 115 230 228 1.1
R62 221 143 1E4
C23 143 115 3.1E-12
C27 227 226 200E-15
C28 225 113 200E-15
R74 4 3 5.0E6
G12 3 4 242 0 -3E-3
I20 0 243 1E-3
D20 243 0 DB
V24 243 194 0.71
R75 0 194 1E6
I21 3 4 115E-6
E25 244 0 120 0 1
C30 114 245 45.0E-12
R78 245 244 25
R81 114 244 1.1E9
I63 0 246 1E-3
D23 246 0 DD
R207 0 246 10E6
V81 246 247 1.798
R208 0 247 2E7
E52 248 0 247 0 -0.875
R209 0 248 1E7
R212 0 247 2E7
G14 237 112 122 0 750E-6
D24 249 250 DL
V42 250 0 3
R213 0 249 3.3E7
G51 2 0 249 0 12.98E-9
I64 2 0 -3.0E-12
G52 212 0 249 0 12.72E-9
I65 212 0 -5.0E-12
G56 118 119 122 0 250E-6
R245 0 120 1E9
S1 120 3 120 3 VSWC
S2 114 110 114 110 VSWC
S3 112 114 112 114 VSWC
S4 251 115 251 115 VSWC
S5 115 252 115 252 VSWC
S6 4 120 4 120 VSWC
E68 116 115 VALUE = {LIMIT(V(114,115),-100,0)}
E69 117 115 VALUE = {LIMIT(V(114,115),0,100)}
R255 115 116 1E9
R256 115 117 1E9
E70 110 111 VALUE = {V(115,116)-V(118,110)}
R157 111 110 1E9
E71 232 112 VALUE = {V(117,115)-V(112,119)}
R158 112 232 1E9
E72 200 112 204 112 50
E73 202 110 203 110 50
V59 253 112 0.30
V60 110 254 1.65
V61 110 238 -1.85
E89 129 0 110 112 1
R203 0 129 1E7
R210 115 144 1E12
G58 3 4 122 0 530E-16
V70 122 0 1
E92 255 256 257 0 1.12E-3
V71 247 257 -1
E93 209 255 258 0 -1.2E-7
R113 0 258 1E9
D25 239 198 DB
R217 0 257 1E12
R220 0 258 1E9
R230 V1 110 1E3
R231 259 V1 60E3
R232 V2 259 60E3
R233 112 V2 1E3
E97 VB1 0 VALUE = {LIMIT(V(VC2),V(VC3),99)}
R234 0 VB1 1E9
E98 VB2 0 VALUE = {LIMIT(V(VC1),-99,V(VC3))}
R235 0 VB2 1E9
E99 VC1 0 VALUE = {4*(V(V1A)-V(VCM))}
R236 0 VC1 1E9
E100 VC2 0 VALUE = {4*(V(V2A)-V(VCM))}
R237 0 VC2 1E9
E101 VC3 0 VALUE = {V(VCM)*(-1)*0.25}
R238 0 VC3 1E9
E102 VB3 0 VALUE = {LIMIT(V(VC3),V(VB2),V(VB1))}
R239 0 VB3 1E9
E103 COUT 0 VALUE = {V(VB1)+V(VB2)}
R240 0 COUT 1E9
E104 V1A 0 VALUE = {(0.75+0.125)*V(V1)}
R241 0 V1A 1E9
E105 V2A 0 VALUE = {(0.75+0.125)*V(V2)}
R242 0 V2A 1E9
S8 220 0 220 0 VSWI
S9 0 220 0 220 VSWI
R246 207 213 100
R247 0 213 1E12
R248 208 214 100
R249 0 214 1E12
E106 242 0 VALUE = {V(194)*0.3+ (V(4)-V(3))*(V(4)-V(3))*(-7E-6)}
R250 0 242 1E9
V79 251 114 -1.2
V80 114 252 -1.2
E109 254 240 194 0 1.25
E110 241 253 194 0 1.25
S10 230 228 260 231 VSWV
S11 230 228 231 261 VSWV
S12 230 228 260 212 VSWV
S13 230 228 212 261 VSWV
V82 110 260 1.25
R156 260 110 1E12
V83 261 112 -0.1
R257 112 261 1E12
R258 120 5 0.1
E111 233 115 VALUE = {LIMIT(V(143,115),V(STN)*0.95,V(STP)*0.85)}
R259 115 233 1E9
R159 212 262 413
R160 262 235 413
C31 262 0 1.2E-14
R161 263 256 413
R162 231 263 413
C32 263 0 1.2E-14
G59 3 4 3 4 -2.0E-6
E113 258 0 VALUE = {(12/(V(VCK))*V(COUT))}
R277 0 258 1E9
E114 VCL 0 VALUE = {LIMIT((SQRT(V(3)-V(4))+1),2.68,6.30)}
R278 0 VCL 1E9
E116 VCK 0 VALUE = {V(VCL)*3-8.5}
R280 0 VCK 1E9
E117 STP 0 VALUE = {((V(194)+0.044)*(-0.4))+0.383}
R284 0 STP 1E9
E118 0 STN VALUE = {((V(194)+0.044)*(-0.4))+0.383}
R285 STN 0 1E9
I11 0 211 0.2E-6
I10 0 210 0.2E-6
D9 210 0 DVN
D10 211 0 DVN
D26 229 264 DIZ
D27 231 264 DIZ
.MODEL NOUT NMOS (LEVEL=3 PHI=0.7 TOX=2E-8 XJ=5E-7
+ TPG=1 VTO=0.5 DELTA=0.5 LD=1E-7 KP=2E-4 UO=650
+ THETA=0.1 GAMMA=0.5 NSUB=1E17 NFS=6E11 FC=0.5
+ VMAX=1E5 ETA=3E-6 KAPPA=10 PB=1 IS=1E-18)
.MODEL POUT PMOS (LEVEL=3 PHI=0.7 TOX=2E-8 XJ=5E-7
+ TPG=-1 VTO=-0.5 DELTA=0.5 LD=1E-7 KP=2E-4 UO=650
+ THETA=0.1 GAMMA=0.5 NSUB=1E17 NFS=6E11 FC=0.5
+ VMAX=1E5 ETA=3E-6 KAPPA=10 PB=1 IS=1E-18)
.MODEL DVN D KF=1.45E-14 IS=1E-16 RS=2E6
.MODEL DIN D KF=3E-15 IS=1E-16 RS=949E3
.MODEL DIZ D IS=1E-18 RS=174
.MODEL PIN PMOS KP=200U VTO=-0.7
.MODEL NIN NMOS KP=200U VTO=0.7
.MODEL HVP PMOS KP=200U VTO=-0.7
.MODEL DL D IS=0.95E-12 N=1.47 XTI=3.5
.MODEL DD D CJO=0.1E-12 TT=10E-9 RS=10
.MODEL DB D CJO=0.1E-12 TT=10E-9 RS=10
.MODEL JC NJF VTO=-0.7 BETA=1E-4 CGS=0.03E-12
+ CGD=0.03E-12 RD=10 RS=10 IS=1E-18
.MODEL QN NPN
.MODEL QP PNP
.MODEL VSWV VSWITCH VON=-0.05 VOFF=0.05 RON=1E-3 ROFF=1E8
.MODEL VSWC VSWITCH VON=0.71 VOFF=0.62 RON=10 ROFF=1E12
.MODEL VSWI VSWITCH VON=0.11 VOFF=0.02 RON=1 ROFF=1E11
.ENDS
* END MODEL NCS2007
